library verilog;
use verilog.vl_types.all;
entity loadarbitrator_demux_sv_unit is
end loadarbitrator_demux_sv_unit;
