library verilog;
use verilog.vl_types.all;
entity shf_sv_unit is
end shf_sv_unit;
