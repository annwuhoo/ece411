library verilog;
use verilog.vl_types.all;
entity comparator_v_sv_unit is
end comparator_v_sv_unit;
