library verilog;
use verilog.vl_types.all;
entity checklruway_sv_unit is
end checklruway_sv_unit;
