library verilog;
use verilog.vl_types.all;
entity lru_way_arbitrator_sv_unit is
end lru_way_arbitrator_sv_unit;
