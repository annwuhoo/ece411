library verilog;
use verilog.vl_types.all;
entity lineoverwrite_sv_unit is
end lineoverwrite_sv_unit;
