library verilog;
use verilog.vl_types.all;
entity lshf_sv_unit is
end lshf_sv_unit;
