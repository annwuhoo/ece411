library verilog;
use verilog.vl_types.all;
entity rshfa_sv_unit is
end rshfa_sv_unit;
