library verilog;
use verilog.vl_types.all;
entity array8_sv_unit is
end array8_sv_unit;
