library verilog;
use verilog.vl_types.all;
entity linetruncate_sv_unit is
end linetruncate_sv_unit;
