library verilog;
use verilog.vl_types.all;
entity shf is
    port(
        \in\            : in     vl_logic_vector(15 downto 0);
        imm4            : in     vl_logic_vector(3 downto 0);
        dbit            : in     vl_logic;
        abit            : in     vl_logic;
        \out\           : out    vl_logic_vector(15 downto 0)
    );
end shf;
