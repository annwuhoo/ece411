library verilog;
use verilog.vl_types.all;
entity cachehit_decoder_sv_unit is
end cachehit_decoder_sv_unit;
