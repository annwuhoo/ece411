library verilog;
use verilog.vl_types.all;
entity pmemconstruct_sv_unit is
end pmemconstruct_sv_unit;
