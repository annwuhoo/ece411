library verilog;
use verilog.vl_types.all;
entity rshfl_sv_unit is
end rshfl_sv_unit;
