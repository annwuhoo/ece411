library verilog;
use verilog.vl_types.all;
entity clonelowbyte_sv_unit is
end clonelowbyte_sv_unit;
