import lc3b_types::*;

module cache_controller
(
    input clk,

	
);



endmodule : cache_controller